module uvm_sepuence_item () endmodule
